interface CpuInterface;
    
endinterface //CpuInterface